askjdasodshadkajhdkjdafdsfsfds