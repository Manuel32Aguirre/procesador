library verilog;
use verilog.vl_types.all;
entity procesador_vlg_vec_tst is
end procesador_vlg_vec_tst;
