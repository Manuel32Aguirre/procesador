LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY dec5_32 IS
	PORT(sel_w_d: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			en_w:IN STD_LOGIC;
			O: OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
END dec5_32;

ARCHITECTURE behavioral OF dec5_32 IS
BEGIN
	PROCESS(sel_w_d)
	BEGIN	
	IF(en_w='1') THEN
	CASE sel_w_d IS
		WHEN "00000" => O <= X"00000001";
		WHEN "00001" => O <= X"00000002";
		WHEN "00010" => O <= X"00000004";
		WHEN "00011" => O <= X"00000008";
		WHEN "00100" => O <= X"00000010";
		WHEN "00101" => O <= X"00000020";
		WHEN "00110" => O <= X"00000040";
		WHEN "00111" => O <= X"00000080";
		WHEN "01000" => O <= X"00000100";
		WHEN "01001" => O <= X"00000200";
		WHEN "01010" => O <= X"00000400";
		WHEN "01011" => O <= X"00000800";
		WHEN "01100" => O <= X"00001000";
		WHEN "01101" => O <= X"00002000";
		WHEN "01110" => O <= X"00004000";
		WHEN "01111" => O <= X"00008000";
		WHEN "10000" => O <= X"00010000";
		WHEN "10001" => O <= X"00020000";
		WHEN "10010" => O <= X"00040000";
		WHEN "10011" => O <= X"00080000";
		WHEN "10100" => O <= X"00100000";
		WHEN "10101" => O <= X"00200000";
		WHEN "10110" => O <= X"00400000";
		WHEN "10111" => O <= X"00800000";
		WHEN "11000" => O <= X"01000000";
		WHEN "11001" => O <= X"02000000";
		WHEN "11010" => O <= X"04000000";
		WHEN "11011" => O <= X"08000000";
		WHEN "11100" => O <= X"10000000";
		WHEN "11101" => O <= X"20000000";
		WHEN "11110" => O <= X"40000000";
		WHEN OTHERS  => O	<= X"80000000";
	END CASE;
	ELSE
	O<=X"00000000";
	END IF;
	END PROCESS;
END behavioral;
		
		
	