averaverque paso aqui