askjdasodshadkajhdkj